.title KiCad schematic
Q1 c b 0 2n2222
V1 bb 0 1v
V2 c 0 10
R1 b bb 1k
.model 2N2222 NPN( Vtf=1.7 Cjc=7.306p Nc=2 Tr=46.91n Ne=1.307
+ Cje=22.01p Vjc=.75 Xtb=1.5 Rb=10 Rc=1
+ Tf=411.1p Xti=3 Ikr=0 Bf=400 Fc=.5
+ Ikf=.2847 Br=6.092 Mje=.377 Mjc=.3416 Vaf=74.03
+ Isc=0 Ise=14.34f Xtf=3 Vje=.75 Is=14.34f
+ Itf=.6 Eg=1.14 )
.dc V2 0 10 0.1 V2 0 10 1
.control
run
plot -i(v2)
.endc
.end
